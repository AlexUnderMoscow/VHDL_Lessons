
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
entity sinlut is
    Port ( en : in  STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (9 downto 0);
           sin : out  STD_LOGIC_VECTOR (11 downto 0));
end sinlut;

architecture Behavioral of sinlut is
type rom_type is array (0 to 1023) of std_logic_vector(11 downto 0);
constant rom: rom_type:=(
x"000",
x"00c",
x"019",
x"025",
x"032",
x"03e",
x"04b",
x"057",
x"064",
x"070",
x"07d",
x"08a",
x"096",
x"0a3",
x"0af",
x"0bc",
x"0c8",
x"0d5",
x"0e1",
x"0ee",
x"0fa",
x"107",
x"113",
x"11f",
x"12c",
x"138",
x"145",
x"151",
x"15d",
x"16a",
x"176",
x"183",
x"18f",
x"19b",
x"1a7",
x"1b4",
x"1c0",
x"1cc",
x"1d8",
x"1e5",
x"1f1",
x"1fd",
x"209",
x"215",
x"221",
x"22e",
x"23a",
x"246",
x"252",
x"25e",
x"26a",
x"276",
x"282",
x"28e",
x"299",
x"2a5",
x"2b1",
x"2bd",
x"2c9",
x"2d4",
x"2e0",
x"2ec",
x"2f8",
x"303",
x"30f",
x"31a",
x"326",
x"332",
x"33d",
x"348",
x"354",
x"35f",
x"36b",
x"376",
x"381",
x"38d",
x"398",
x"3a3",
x"3ae",
x"3b9",
x"3c4",
x"3d0",
x"3db",
x"3e6",
x"3f0",
x"3fb",
x"406",
x"411",
x"41c",
x"427",
x"431",
x"43c",
x"447",
x"451",
x"45c",
x"466",
x"471",
x"47b",
x"486",
x"490",
x"49a",
x"4a4",
x"4af",
x"4b9",
x"4c3",
x"4cd",
x"4d7",
x"4e1",
x"4eb",
x"4f5",
x"4ff",
x"508",
x"512",
x"51c",
x"525",
x"52f",
x"539",
x"542",
x"54b",
x"555",
x"55e",
x"567",
x"571",
x"57a",
x"583",
x"58c",
x"595",
x"59e",
x"5a7",
x"5b0",
x"5b9",
x"5c1",
x"5ca",
x"5d3",
x"5db",
x"5e4",
x"5ec",
x"5f5",
x"5fd",
x"605",
x"60e",
x"616",
x"61e",
x"626",
x"62e",
x"636",
x"63e",
x"645",
x"64d",
x"655",
x"65d",
x"664",
x"66c",
x"673",
x"67b",
x"682",
x"689",
x"690",
x"697",
x"69f",
x"6a6",
x"6ac",
x"6b3",
x"6ba",
x"6c1",
x"6c8",
x"6ce",
x"6d5",
x"6db",
x"6e2",
x"6e8",
x"6ee",
x"6f5",
x"6fb",
x"701",
x"707",
x"70d",
x"713",
x"718",
x"71e",
x"724",
x"72a",
x"72f",
x"735",
x"73a",
x"73f",
x"745",
x"74a",
x"74f",
x"754",
x"759",
x"75e",
x"763",
x"767",
x"76c",
x"771",
x"775",
x"77a",
x"77e",
x"783",
x"787",
x"78b",
x"78f",
x"793",
x"797",
x"79b",
x"79f",
x"7a3",
x"7a6",
x"7aa",
x"7ae",
x"7b1",
x"7b4",
x"7b8",
x"7bb",
x"7be",
x"7c1",
x"7c4",
x"7c7",
x"7ca",
x"7cd",
x"7cf",
x"7d2",
x"7d5",
x"7d7",
x"7da",
x"7dc",
x"7de",
x"7e0",
x"7e2",
x"7e5",
x"7e6",
x"7e8",
x"7ea",
x"7ec",
x"7ee",
x"7ef",
x"7f1",
x"7f2",
x"7f3",
x"7f5",
x"7f6",
x"7f7",
x"7f8",
x"7f9",
x"7fa",
x"7fb",
x"7fb",
x"7fc",
x"7fd",
x"7fd",
x"7fe",
x"7fe",
x"7fe",
x"7fe",
x"7fe",
x"7ff",
x"7fe",
x"7fe",
x"7fe",
x"7fe",
x"7fe",
x"7fd",
x"7fd",
x"7fc",
x"7fb",
x"7fb",
x"7fa",
x"7f9",
x"7f8",
x"7f7",
x"7f6",
x"7f5",
x"7f3",
x"7f2",
x"7f1",
x"7ef",
x"7ee",
x"7ec",
x"7ea",
x"7e8",
x"7e6",
x"7e5",
x"7e2",
x"7e0",
x"7de",
x"7dc",
x"7da",
x"7d7",
x"7d5",
x"7d2",
x"7cf",
x"7cd",
x"7ca",
x"7c7",
x"7c4",
x"7c1",
x"7be",
x"7bb",
x"7b8",
x"7b4",
x"7b1",
x"7ae",
x"7aa",
x"7a6",
x"7a3",
x"79f",
x"79b",
x"797",
x"793",
x"78f",
x"78b",
x"787",
x"783",
x"77e",
x"77a",
x"775",
x"771",
x"76c",
x"767",
x"763",
x"75e",
x"759",
x"754",
x"74f",
x"74a",
x"745",
x"73f",
x"73a",
x"735",
x"72f",
x"72a",
x"724",
x"71e",
x"718",
x"713",
x"70d",
x"707",
x"701",
x"6fb",
x"6f5",
x"6ee",
x"6e8",
x"6e2",
x"6db",
x"6d5",
x"6ce",
x"6c8",
x"6c1",
x"6ba",
x"6b3",
x"6ac",
x"6a6",
x"69f",
x"697",
x"690",
x"689",
x"682",
x"67b",
x"673",
x"66c",
x"664",
x"65d",
x"655",
x"64d",
x"645",
x"63e",
x"636",
x"62e",
x"626",
x"61e",
x"616",
x"60e",
x"605",
x"5fd",
x"5f5",
x"5ec",
x"5e4",
x"5db",
x"5d3",
x"5ca",
x"5c1",
x"5b9",
x"5b0",
x"5a7",
x"59e",
x"595",
x"58c",
x"583",
x"57a",
x"571",
x"567",
x"55e",
x"555",
x"54b",
x"542",
x"539",
x"52f",
x"525",
x"51c",
x"512",
x"508",
x"4ff",
x"4f5",
x"4eb",
x"4e1",
x"4d7",
x"4cd",
x"4c3",
x"4b9",
x"4af",
x"4a4",
x"49a",
x"490",
x"486",
x"47b",
x"471",
x"466",
x"45c",
x"451",
x"447",
x"43c",
x"431",
x"427",
x"41c",
x"411",
x"406",
x"3fb",
x"3f0",
x"3e6",
x"3db",
x"3d0",
x"3c4",
x"3b9",
x"3ae",
x"3a3",
x"398",
x"38d",
x"381",
x"376",
x"36b",
x"35f",
x"354",
x"349",
x"33d",
x"332",
x"326",
x"31a",
x"30f",
x"303",
x"2f8",
x"2ec",
x"2e0",
x"2d4",
x"2c9",
x"2bd",
x"2b1",
x"2a5",
x"299",
x"28e",
x"282",
x"276",
x"26a",
x"25e",
x"252",
x"246",
x"23a",
x"22e",
x"221",
x"215",
x"209",
x"1fd",
x"1f1",
x"1e5",
x"1d8",
x"1cc",
x"1c0",
x"1b4",
x"1a7",
x"19b",
x"18f",
x"183",
x"176",
x"16a",
x"15d",
x"151",
x"145",
x"138",
x"12c",
x"11f",
x"113",
x"107",
x"0fa",
x"0ee",
x"0e1",
x"0d5",
x"0c8",
x"0bc",
x"0af",
x"0a3",
x"096",
x"08a",
x"07d",
x"070",
x"064",
x"057",
x"04b",
x"03e",
x"032",
x"025",
x"019",
x"00c",
x"000",
x"ff4",
x"fe7",
x"fdb",
x"fce",
x"fc2",
x"fb5",
x"fa9",
x"f9c",
x"f90",
x"f83",
x"f76",
x"f6a",
x"f5d",
x"f51",
x"f44",
x"f38",
x"f2b",
x"f1f",
x"f12",
x"f06",
x"ef9",
x"eed",
x"ee1",
x"ed4",
x"ec8",
x"ebb",
x"eaf",
x"ea3",
x"e96",
x"e8a",
x"e7d",
x"e71",
x"e65",
x"e59",
x"e4c",
x"e40",
x"e34",
x"e28",
x"e1b",
x"e0f",
x"e03",
x"df7",
x"deb",
x"ddf",
x"dd2",
x"dc6",
x"dba",
x"dae",
x"da2",
x"d96",
x"d8a",
x"d7e",
x"d72",
x"d67",
x"d5b",
x"d4f",
x"d43",
x"d37",
x"d2c",
x"d20",
x"d14",
x"d08",
x"cfd",
x"cf1",
x"ce6",
x"cda",
x"cce",
x"cc3",
x"cb8",
x"cac",
x"ca1",
x"c95",
x"c8a",
x"c7f",
x"c73",
x"c68",
x"c5d",
x"c52",
x"c47",
x"c3c",
x"c30",
x"c25",
x"c1a",
x"c10",
x"c05",
x"bfa",
x"bef",
x"be4",
x"bd9",
x"bcf",
x"bc4",
x"bb9",
x"baf",
x"ba4",
x"b9a",
x"b8f",
x"b85",
x"b7a",
x"b70",
x"b66",
x"b5c",
x"b51",
x"b47",
x"b3d",
x"b33",
x"b29",
x"b1f",
x"b15",
x"b0b",
x"b01",
x"af8",
x"aee",
x"ae4",
x"adb",
x"ad1",
x"ac7",
x"abe",
x"ab5",
x"aab",
x"aa2",
x"a99",
x"a8f",
x"a86",
x"a7d",
x"a74",
x"a6b",
x"a62",
x"a59",
x"a50",
x"a47",
x"a3f",
x"a36",
x"a2d",
x"a25",
x"a1c",
x"a14",
x"a0b",
x"a03",
x"9fb",
x"9f2",
x"9ea",
x"9e2",
x"9da",
x"9d2",
x"9ca",
x"9c2",
x"9bb",
x"9b3",
x"9ab",
x"9a3",
x"99c",
x"994",
x"98d",
x"985",
x"97e",
x"977",
x"970",
x"969",
x"961",
x"95a",
x"954",
x"94d",
x"946",
x"93f",
x"938",
x"932",
x"92b",
x"925",
x"91e",
x"918",
x"912",
x"90b",
x"905",
x"8ff",
x"8f9",
x"8f3",
x"8ed",
x"8e8",
x"8e2",
x"8dc",
x"8d6",
x"8d1",
x"8cb",
x"8c6",
x"8c1",
x"8bb",
x"8b6",
x"8b1",
x"8ac",
x"8a7",
x"8a2",
x"89d",
x"899",
x"894",
x"88f",
x"88b",
x"886",
x"882",
x"87d",
x"879",
x"875",
x"871",
x"86d",
x"869",
x"865",
x"861",
x"85d",
x"85a",
x"856",
x"853",
x"84f",
x"84c",
x"848",
x"845",
x"842",
x"83f",
x"83c",
x"839",
x"836",
x"833",
x"831",
x"82e",
x"82b",
x"829",
x"826",
x"824",
x"822",
x"820",
x"81e",
x"81b",
x"81a",
x"818",
x"816",
x"814",
x"812",
x"811",
x"80f",
x"80e",
x"80d",
x"80b",
x"80a",
x"809",
x"808",
x"807",
x"806",
x"805",
x"805",
x"804",
x"803",
x"803",
x"802",
x"802",
x"802",
x"802",
x"802",
x"801",
x"802",
x"802",
x"802",
x"802",
x"802",
x"803",
x"803",
x"804",
x"805",
x"805",
x"806",
x"807",
x"808",
x"809",
x"80a",
x"80b",
x"80d",
x"80e",
x"80f",
x"811",
x"812",
x"814",
x"816",
x"818",
x"81a",
x"81b",
x"81e",
x"820",
x"822",
x"824",
x"826",
x"829",
x"82b",
x"82e",
x"831",
x"833",
x"836",
x"839",
x"83c",
x"83f",
x"842",
x"845",
x"848",
x"84c",
x"84f",
x"852",
x"856",
x"85a",
x"85d",
x"861",
x"865",
x"869",
x"86d",
x"871",
x"875",
x"879",
x"87d",
x"882",
x"886",
x"88b",
x"88f",
x"894",
x"899",
x"89d",
x"8a2",
x"8a7",
x"8ac",
x"8b1",
x"8b6",
x"8bb",
x"8c1",
x"8c6",
x"8cb",
x"8d1",
x"8d6",
x"8dc",
x"8e2",
x"8e7",
x"8ed",
x"8f3",
x"8f9",
x"8ff",
x"905",
x"90b",
x"912",
x"918",
x"91e",
x"925",
x"92b",
x"932",
x"938",
x"93f",
x"946",
x"94d",
x"954",
x"95a",
x"961",
x"969",
x"970",
x"977",
x"97e",
x"985",
x"98d",
x"994",
x"99c",
x"9a3",
x"9ab",
x"9b3",
x"9bb",
x"9c2",
x"9ca",
x"9d2",
x"9da",
x"9e2",
x"9ea",
x"9f2",
x"9fb",
x"a03",
x"a0b",
x"a14",
x"a1c",
x"a25",
x"a2d",
x"a36",
x"a3f",
x"a47",
x"a50",
x"a59",
x"a62",
x"a6b",
x"a74",
x"a7d",
x"a86",
x"a8f",
x"a99",
x"aa2",
x"aab",
x"ab5",
x"abe",
x"ac7",
x"ad1",
x"adb",
x"ae4",
x"aee",
x"af8",
x"b01",
x"b0b",
x"b15",
x"b1f",
x"b29",
x"b33",
x"b3d",
x"b47",
x"b51",
x"b5c",
x"b66",
x"b70",
x"b7a",
x"b85",
x"b8f",
x"b9a",
x"ba4",
x"baf",
x"bb9",
x"bc4",
x"bcf",
x"bd9",
x"be4",
x"bef",
x"bfa",
x"c05",
x"c10",
x"c1a",
x"c25",
x"c30",
x"c3c",
x"c47",
x"c52",
x"c5d",
x"c68",
x"c73",
x"c7f",
x"c8a",
x"c95",
x"ca1",
x"cac",
x"cb7",
x"cc3",
x"cce",
x"cda",
x"ce6",
x"cf1",
x"cfd",
x"d08",
x"d14",
x"d20",
x"d2c",
x"d37",
x"d43",
x"d4f",
x"d5b",
x"d67",
x"d72",
x"d7e",
x"d8a",
x"d96",
x"da2",
x"dae",
x"dba",
x"dc6",
x"dd2",
x"ddf",
x"deb",
x"df7",
x"e03",
x"e0f",
x"e1b",
x"e28",
x"e34",
x"e40",
x"e4c",
x"e59",
x"e65",
x"e71",
x"e7d",
x"e8a",
x"e96",
x"ea3",
x"eaf",
x"ebb",
x"ec8",
x"ed4",
x"ee1",
x"eed",
x"ef9",
x"f06",
x"f12",
x"f1f",
x"f2b",
x"f38",
x"f44",
x"f51",
x"f5d",
x"f6a",
x"f76",
x"f83",
x"f90",
x"f9c",
x"fa9",
x"fb5",
x"fc2",
x"fce",
x"fdb",
x"fe7",
x"ff4"
);
begin
rom_select: process (addr,en)
begin
	if (en='0') then
		sin <= "000000000000";
	else
		sin <= rom(conv_integer(addr));
	end if;
end process;
end Behavioral;

